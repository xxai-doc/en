�TV����.h�����,�\�	��96���